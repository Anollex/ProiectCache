library verilog;
use verilog.vl_types.all;
entity controlUnitCache_tb is
end controlUnitCache_tb;
